----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/30/2019 02:26:36 AM
-- Design Name: 
-- Module Name: 4BitRegister - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FourBitRegister is
    Port ( D : in STD_LOGIC_VECTOR (3 downto 0);
           Load : in STD_LOGIC;
           clr : in STD_LOGIC;
           clk : in STD_LOGIC;
           Q : out STD_LOGIC_VECTOR (3 downto 0));
end FourBitRegister;

architecture Behavioral of FourBitRegister is

begin

process (clk, D) is
    begin
        if (clk'event and clk ='1') then
            if (clr ='1') then
                Q <= (others => '0');
            elsif (Load = '1') then
                Q <= D;
            end if;
        end if;
    end process;

end Behavioral;
